`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
//Students: Brett Bushnell (Undergrad), Matt Dzurick (Grad)
//Date Created: Mon Oct 24 20:07:17 2016


//Assignment: 2
//File: 474a_circuit1_output.v
//Description: Netlist Behavior circuit implementation for C:\Users\Brett\Dropbox\School_F2016\ECE474A\Assignment2\assignment_2_circuits\474a_circuit1_output.v
//
//////////////////////////////////////////////////////////////////////////////////


module 474a_circuit1_output(Clk, Rst, a, b, cz, x);
	input [7:0] a;
	input [7:0] b;
	input [7:0] c;

	output [7:0] z;
	output [15:0] x;

	wire [7:0] d;
	wire [7:0] e;
	wire [15:0] f;
	wire [15:0] g;
	wire [15:0] xwire;


endmodule
